module IDEX_
